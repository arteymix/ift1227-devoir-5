library ieee; use ieee.std_logic_1164.all;

entity snail is
    port(
        clk:    in std_logic;
        input:  in std_logic;
        output: out std_logic
    );
end entity;

architecture sticky of snail is
begin

    

end architecture;
